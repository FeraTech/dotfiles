BSV1    �`y��U  FCS��U  U&      H  PC     [�A      �X      Y      &S      �P      �DB     �RAM    �HJ �     -  �Ɍ97E+���X    diTJ                                      (	  �  ��  &2� �wL ��j"`�Pp�&%� M:�` A0��mm�c���mm� ���� ��    �                    �                                        � dd� ��� Z       ������������� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������N�~~�7�4�}�x�x��r�[��a X�  �  �  �  �  �  ���B��  �  �  �  �  �  �  ��d���� ��T ��> �/> !�>2��h����c�¨��Ahm�*m�r��B�H��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �m�jm�"��A`c����� ��� �6������ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �? �����efff$ ��������� l! �!$ �!$�                     x� �N͉    		                                                             �� �               @ ��               `@ @ @   ���                                                             p�p�p                   �����                                                            o.                       ������&&&&&&&&&��&                         ���                                                                                       ��Z      ������������������������������������������������                                                                                                                                                ��� �                  G��L		0		 (  STdD4R         �    


$$$$$$$$$$$$$$$$$$$$$��            0�|            �              7    �        �  ���        � �   ���   �!� 00�&  %�"00�0�  �0 �2�p���� $�!����2�:� �0��)*����0� �� 0 �� ��6840 �1����� 0�������a���!�0!2�!��&� $����� �(�0 ��"��  00        �����          �����           4��0            ���             4�0             8��             ������          �       �F   JAMM    IQLB       ICoa       ICou   ����TSBS   A jn   MooP   ��	  NTAR   $$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$��������$�!iki
k$$bb$$$$$��������$$$$$l$ll$l$$$$$$$$$$$$$��������$�!$l$ll$l$���efff$$$$$��������$a!$njmnjm$��������$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$������&&&&��������&&&&����&&����������&&&&��������&&&&����&&����������&&&&��������&&&&����&&����������&&&&����$$��&&&&����&&����������&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&��������������������������������������������������������������������������������������������������������������������������������  @  DUU    DUU������������������������������������������������������&&&&��������&&&&����&&����������&&&&��������&&&&����&&����������&&&&��������&&&&����&&����������&&&&����$$��&&&&����&&����������&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&��&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&������&&&&&&&&&&&&&&&&&&&&&&&&&&��������������������������������������������������������������������������������������������������������������������������������$$$$$$$$$$$$$$$��$$$$$$$$$$$$$$$$$$$$$$$$$$$$$����$$$$$$$$$$$$$$$$$$$$$$$$$$$������$$$$$$$$$$$$$$$$$$$$$$$$$��������$$$$$$$$$$$$$$$$$$$$$$$������$���$$$$$$$$$$$$$$$$$$$$$������������$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$������������������������������������������������UUUUUUUUUUUUUUU�PRAM    0 '677 2' "0 '0 SPRA   �a X�  �  �  �  �  �  ���B��  �  �  �  �  �  �  ��d���� ��T ��> �/> !�>2��hd�����A`m�#m�j���6��H��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �m�rm�+��Ahd�¨�� ��� �H���B��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �PPUR   �  KOOK   DEAD    PSPL    XOFF    VTGL    RADD    TADD     VBUF   �PGEN   �   JYRB    JOYS       LSTS    $  FHCN   �! FCNT    PSG    ���w � ENCH   IQFM   NREG   &@TRIM    TRIC    E0SP   E1SP   E2SP   E0MO   E1MO   E2MO   E0D1   E1D1   E2D1   E0DV   E1DV   E2DV   LEN0   �   LEN1   �   LEN2   �   LEN3       SWEE     CRF1   �   CRF2   w   SWCT   SIRQ    5ACC   6   5BIT   5ADD   }G  5SIZ   d   5SHF   5VDM   5VSP   5SZL   
5ADL   5FMT   RWDA   .SAC1   X8� SAC2   b�RCD1      RCD2      TRIS      TACC   6@ NACC   F�' CBC1      CBC2      CBC3      CBC4      CBC5      SNTS       TSOF      WLC1      WLC2      WLC3      WLC4      FAC1   ��>%    FAC2   G������TCOU       WAVE�                                                                                                                                 >@  CHRR     w�9   	>>~��p ??��p ����    ������44t���p��ܔ$�pw�9  	 ?xxy? w~ ����"" ������������� �>"�  �

 9  '/=??7# ����PP�  ������>�����p ���� p     0<??00 ��������  <x�������` � `  8|N   ?��p ��p ������   x������������|����/o��j98s���w3;  8  ����xX��  �����<���� �<�p��� ?__@``pxmg???��    O��  ��������   8�ӿ������<<??>�<<                                ���                  ���        88888888888888888��8 8888 8 8 ,<~��, T�_�V<4�( 4  <tn$ <<   <<<<<<<<  <=====�~       ***  """������������������ �(.|�x        xxB����8|Ƃ���Hpp0p   x����   x������`p0   ��pp0   0p�����<~���������   �����~<<N 0����~<  p`          80    Pp    pp8        @@`�    ���H     8|?          �B      ���`      ?<         D-�|    D-�|8|�    8|�    ���                              <<$$f�< <$$$f��������~�������~�������� �������������~�����      <~f��     <<��f~<   <<        >>      A>A       `Ab<    ����pp4:����pp0:_N, H<<<    $           5+^�������<|X�����x�� :s�1� t���0�pq �� 
2 8T���nF(D(���R:T8|    l�*80   8T~FG�ǮD( 8y���9    F�(80   ����#" ��������������?#��  ���灁  ����������~<  ����~<  

   '/=?|ߍ��������~

 	  '/=?>oFnn~  ?>  )+-{z    Br���ss< D�������       �_F���@������ 

��  '/=?��灁���~<������~<   
   
      @ �@!	�� @�	!@?   ?/??   >>?  "A@@@?       	''#  8?;18?       1{{{{{1{{{@;{{{{{{N  {{@;{{{1                      ?woo��?����[��??)#0v�+#0v��)#k1
�k#k1
   
   
�	  �	   �������������������������������ojb09=`sg}??; ?p@�       <     `@     �@` 0  0 `@�    ����`` ``����   ����&$  ������44t���v��ޖ&�v     �       W��    WW             �       ���      ��           �T�     �T T�      T�             �                                    �        �             _      �_      �      ?ww~����������������om}}��������>	 %>~11qa ^^^^, � 88 �������������`X|x��`     p C  ��S0  >6
 � 0� >4 �0 �0 ���<���  
  <www/���    8< 
~^__Wo/!	)   $??/gOGppya  d���  8|����N~    ��~    	��������������� ������ ���
��uu��
���~�&�8�>��>	��������������� ������  ���
��uw��
���{�& �;�>��<���@O`(���O@__( ?@@`D@_���?_x@H(00?�{9�������=?�???����� p���D@O (���OO@__( @@@|�߀_@8H(00?�{9�������=?�?? ���Ɔp �}7�? _	     �o=�?�3  	      ����    ����     $l������   ��"H�������l$�H"��   	'7??    ??7'	    �������   ��"H���������H"��                              7                                        �=/;^wP!!#7?! 19	7=o��		A" }�}#~�c!0    8}?< 8|>?<x 0?      ಀ�    �?� ������7?�    h@G W?>�3pB@@@�B    ���?�         ��>?>  xp����������      �    �   ��??       �xP@>?  ������>��������       
4{���|@�	`````@��� �@����\�`�����xp�,   	  {��=??? �l     �����@   �����x���xpX@�         ?7    <~��7?    ��~    ����c����\  ???   ��b������x�~��x0��������0����>  �oo?�????~��??�  �������������������� ��������    	3#G.\]����@  ��o? �0�����������FLLx��x8����  ���������Aej�jjo�����L#�\X�/#���������Aem�uuu�����O#�um�-!  >?xx  Gqpxy?# >�??  ��������{o�������>>�  |   >?y   xx|~<8 G7 �   � ������{�@ p o������ Wa$'$<N^_\�Px?T��GP;|| (`��&�$<ؠpx�:ڈ���� v���    '?<( ``@? @@XG <<   �����<��������� 6� 8L���d8         8~         |�<x��         ~<�|         <l��         ����|         <`����|         ��000         x��x��|         |��~x         8l�����         �������         <f���f<         �������         �������         �������         >`���f>         �������         <<         ��|         �������         ``````~         �������         �������         |�����|         �������         |�����z         �������         x��|�|         ~         ������|         ����|8         �������         ��|8|��         fff<         �8p��                         ��������                ������������������������    0                    0              p�P T�v              00         $$$             8D             �            �_UUU   �_UUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   .__�~< <^���~<   �                 00         �         l����|8 l����|8l����|8���     ���     � B ��������         ��      ��      ��   ����   ��         �� ��� �  ��  ����������  ``nnnn��������nnnnnnn �      ���������� ??????������������������������������       ��������       �������������������     ��������        ��������        ���������O��������      ��������       �����������������O���        ��������        ��������       ���������������    @ ��������    � �����}��  @  ��������    @���������������������o���3�YBR���?������������������������mIN�ok;o���������~����������   ��������?۟������  c������ c��������������������  ��������������������~�������������������? �������������������������������������o������������������������ �����s��  ������ ������ �����hh��hh�����x3A�        ��������<~����@ Á�� ?//��������////??��������������������������� ������ � ||8x  �����~������ ������� ����������������������~ ������ ��������  |�  ����0   ?@�� ��������  >@@@���@@ �      ����1     xp�񹩩�                ��������        ��������-----��������iK[[_��̀����  2Fx8~�7��������   ����������������  ����Ǉ     ���  ������      �����䄀          /�       �����>      ��������        ��������        +V�� ���Ç@ ��   @??????3��������������� Ã���   ���px��?��~zz���� 


�   '��������    ������     � �������O�������<| ����  
/7}��������  ���~ �   ����  �������?d���  � �0xY�����ǃ�BBDsss���} ���   �   ����x`��h((���       ��������6~vtt��������  0x�||x||Á�������||�xL�   8||~~|��Á������|~��� �        �����������||x�����������G�      ���������������Ã �������qs���	����A@���,��  @R��������    !�ޜ�    !!! �~O7wwww��������vv664   ��@@@A?�     !!#?        ���� ??�����x`gH�����2>A��  ����-7����   ����mL� |� ������� �������        ?         �������  @� ?��@  �������� @�  @� @  @   @� @��@ ��@ � @� @��@ ��@ �      �      ��      ��      ��      ��      �l����|8                        ��������                ��������`@@����� ���  @ ��� =}�����                       	 P�� �  ��  ��     ���     ��� <B����B<                ������        ��������� ��� ��� ��� WRAM     Z


$$$$$$$$$$$$$$$$$$$$$  ??    [��?                                                                                             �              7    �          ���      �    �   ��   �!� 00�&  %�"00�0�  �0 �2�p���� $�!����2�:� �0��)*����0� �� 0 �� ��6840 �1����� 0�������a���!�0!2�!��&� $����� �(�0 ��"��  00                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �     ZZZ���R/  ���   ��������&&&&&&����������������&&&&&&����������������&&&&&&����������������&&&&&&��������������&&&&&&&&&&������������&&&&&&&&&&������&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&��&&��&&&&��������&&&&��&&��&&&&�������$&&&&&&&&&&&&&&�������$&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&����&&&&&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&��������&&&&&&&&&&&&&&����?  0 '6,,2')')''0�?
*� Bb�؛�>���Ĝ��2�m����'�l���ߞ!�U�*������+�������+,���������+K
������$����+���cs�S���+s��W��S�#��c�Kk�3'�gPPsC�;����_`pp�Cs�cr�  cK����2���r ��

��

2r�csr
rr2
�RBb�?�SC�*bBRc�oo'_k_k'G_OK{kc�[c�_{[koWS_ZDLSwk�k�G�D h�G
�  v~F�Rvj~� �����z[�_j{�^^�""�ws�_fZBjSG[_ BB��� ��  A��eB��  ���!!B Z���P��N�I !!� O  �/�O
C�	!!/G  P��ĪCC���c�iGiiZGcCC��䃃�iiGGGi�DD�Z�bC�N G�M��IH	 ��	
��� !"#$%&'()�+�-./0�23456�8�:
;�=>?88@ABCD�FG�IJ�LM���QR��UV�XYZ��\]����bcd��gh��kl�no�qrstuvvwx? ?Z??????���????????��XؘX� ����?�?�?�                  


         ( D

2�P�d<Zd
P�<   d  
 ��������� � E� �    �   �  ��� �b   @� �E  �     ��      E 	 
  �  �    �K   @ M�I�  H�   " @    ?  0 '6772'"0'0,��WI�i  w* #Iy������*���������������� bH� �H� �H� �H������������������������������������������������������������������������������������������������������������������������������?                    � ��` �$$$$$$$$ �$$$$$$$$ l! $ �! $ �! $���ҭ͠'�m��&���� �W�J���}��}�m���~��~�m���(��l�����o��p� yn��m� Pm�!�d�� �!��
 um� UmLFm��n Pm��X�'LPm�  dm�� � �ʈ�` Un�$��!��$����$�`��� � `�H Ƈ ���p�p�݅���� <� ��h�� ���0����Z`� �+�,�-``�``eeeeB`b
`eeeej`�c`eeee���i������m� �������`�;�� �m�
�;`�`��� ����� ���B 9n�B`�Ai�(�� �A`��Ɏ���)��LI� nn�� nn� ��$� ����`� �
���
�����H)� �8� � hJJJJ��8��� �i�����	�i�������$�� �������ɀ��� �)�e��f��������й`����
��` �
� �p� �� }�n�����@	 �@����� �� ��`��p� � ����O�\�� i� � �F�� ����O�\�� 8�� �� �G�J�%�ELI���� � ����O�\�� i� � �H��� ����O�\�� 8�!� �� �I��`� )o so�`��}���������((��i ��(`��8����������(8(��� ��(`�J����p`I�i` �o���H� �� ��h��}���`���`H���
�p �p �p��
�h���
�� �� �p�`� ������H��h����8���� e� ����8����� `����)��@�^�ހ��P��`������F
�8��	�� `�X������)���赬�)���B�I��� ���5�X� �� �(����������������� <qep�p��JJ <qe���`� � )��)�ȹ  `����赬���[������� ����� ���!��� �m��� q`���j)0JJJJ���kH)



�h)�`���ӕ(����������`������J�(����*L�q����
��`��	�[�"�V�� H)pJJi�T����� h)� �


e m�k�W�>�U� � ��H��	��q9����)��h�Hh�V` Hr�L���(�'��
�
�|�� ��� �� ި�
�����(�|�}`�e � ��`�e���`�e���`�8����`   	
!"#!"!"!""��         ��	� `��k���k�	��)`)2��)��@�� s����0鵘�����r��i8�� p�	�c�p8�p p�	�W�������� s��������������� ����r���rH)�
h)����r��n��j��f�
�W`� �t��`��M��:�����>��u�� �t��m�
yW�����������|��|L�s�W��iL�sL�t� ���k��-��[�����8�����)��W��W�� ���` �t�
� lt��p��	`�o��`���p`�oH)� hJJJJ� `� ��L���
�W� �W����b�%s��hL+���}`� ���`�4�K�I�� 


e )����?����� ��k���� ��������)���
�4`� `=  �  � � �
u� �)���@��`�/�����a��'u���'�/��`� �/`��� Iu������+u����`��٩�`�� �
& 
& )���JJJ�`���������� \`!!dj')+5?ptvvxz~�I���KOOQQ�����������ST���������������������������������		

�UUUUUUUVWW��XXXXXXXXXYYYYZZZZ[[[ \�D�������������������������������̼���������������������������Ƞ���������ɽ�����������������������������������������  ������������������������������������������������������������������rt������          ����     `�d�h�l�p�t�x�|��܄؈ԌА�����������` O��L�w��� ��Oȅ���A��w�C��w� ��H�C�L�D�����
��ue��v�i�� �����)���)���v �y� ���Lyy�Lhx���H��h��I@��I@������ )�� ��) � ��C� � ��� � �e
� � ��D�� 6n��֦` 
 !""&'()+. �<4prt(�<*&$"@J�lBFv,NLjPRf2.h�n�68:<VHx �z|0db �y� ���H� �R�A��w�C��w�Dh������
��xe���x�i������ ��b���� i� �R� �Lhx�l��|�LNx��
���I@�Lhx���`��H����)��A��w�h��p���� ��L6n �y����� � ��L�w -z��) �#���=� �{� �|� �|� �|� )}� _} �z�O���������,� �O`�'������,`�����)@�F�pe���e�`������������� ����������        ���        ���� -z� �K��	�� � ��l==�t���@�n��i�O�S���)���Z�pi���i��	 �}�E�O�S�?�K�V�8�Z�4��)��.���)��
���)���O�U�	�[��v�
��� �` &~��O�JzH)�h)���O�.�� |m�b�Ff���� �'�P�Q�p��8��p�o)��#�o8��o`�8�p��o)�
�o���pо�o)��o ��p�������`�� 
��� ��	�
���p i��� i�� �� �� �y �}�t����%	� �}�P�� ��%	�Z� ���=��%	�L�O�3��4�L@��������� ��LT|������ �����������8����`�	� �����L�}�'�P�
��P�P�
��	���Q ��� �= ���`� ��	�� J�2���� � 
���	�@�W��� ���� �}��	�H� ��h�`� � �	������ � ���0��	�@����p i��� i�� �}� |��%	� &~` @� ��	�� ���W�%}���)�	���LS}���� �}���L�}� �� �0���	� ��� �V��	� �Y��
�� �}��=���O��� ��LT|� �� ����O������ �����L&~��`���� ��)��p i��� iL�}�p i��� iL�{��� �� �8� p�
���8� p�����`� ����%	�j������� �� ������)��������p��p ����F� �.���(�	������� ������)���O���� p��`�� ���)���	@����+�O�3��4�������k���	����@�ө��`�������������������������������                                                                                                                                                                                                                                                               �DREG     LRST   �]     BFFR    BFRS                                                                                                                